// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Sun May 17 21:05:09 2020

// synthesis message_off 10175

`timescale 1ns/1ns

module TM1638_shifter (reset,clock,data_in,data_io,strobe);

    input reset;
    input clock;
    input [7:0] data_in;
    tri0 reset;
    tri0 [7:0] data_in;
    output data_io;
    output strobe;
    reg data_io;
    reg reg_data_io;
    reg strobe;
    reg [8:0] fstate;
    reg [8:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4,state6=5,state7=6,state8=7,state9=8;

    initial
    begin
        reg_data_io <= 1'b0;
    end

    always @(posedge clock or posedge reset)
    begin
        if (reset) begin
            fstate <= state1;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or data_in or reg_data_io)
    begin
        reg_data_io <= 1'b0;
        strobe <= 1'b0;
        data_io <= 1'b0;
        case (fstate)
            state1: begin
                reg_fstate <= state2;

                strobe <= 1'b0;

                reg_data_io <= data_in[0];
            end
            state2: begin
                reg_fstate <= state3;

                reg_data_io <= data_in[1];
            end
            state3: begin
                reg_fstate <= state4;

                reg_data_io <= data_in[2];
            end
            state4: begin
                reg_fstate <= state5;

                reg_data_io <= data_in[3];
            end
            state5: begin
                reg_fstate <= state6;

                reg_data_io <= data_in[4];
            end
            state6: begin
                reg_fstate <= state7;

                reg_data_io <= data_in[5];
            end
            state7: begin
                reg_fstate <= state8;

                reg_data_io <= data_in[6];
            end
            state8: begin
                reg_fstate <= state9;

                strobe <= 1'b1;

                reg_data_io <= data_in[7];
            end
            state9: begin
                reg_fstate <= state9;

                reg_data_io <= 1'b0;
            end
            default: begin
                reg_data_io <= 1'bx;
                strobe <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
        data_io <= reg_data_io;
    end
endmodule // TM1638
